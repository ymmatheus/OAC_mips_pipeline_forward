library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity mux41 is
	port (
		sel			: in  std_logic_vector(1 downto 0);
		A,B,C			: in  std_logic_vector(31 downto 0);
		S				: out std_logic_vector(31 downto 0));
end mux41;

architecture behavioral of mux41 is

begin
	proc_mux: process(A,B,C,sel) 
	begin
      case sel is

			when  "00" => S <= A;
			
			when  "01" => S <= B;
			
			when	"10" => S <= C;
		
			when others => S <= X"00000000";
	  
	  end case;
	end process proc_mux;
end architecture behavioral;







