-- Unidade de Controle MIPS
-- 					Sinais de Controle
-- Execução/ Calculo endereço: RegDst, OpALU1, opALU0, OrigALU
-- Acesso a Memoria: Branch, LeMem, EscreveMem 
-- Escrita do Resultado: EscreveReg, MemtoReg
 
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
