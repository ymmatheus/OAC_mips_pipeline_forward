-- PC MIPS