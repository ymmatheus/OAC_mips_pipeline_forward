-- PC MIPS



